`timescale 1ns/1ps
// (Optional for SV-only tools; Icarus uses `timescale`)
// timeunit 1ns; timeprecision 1ps;